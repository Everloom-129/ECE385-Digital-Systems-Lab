
module lab7_spc (
	clk_clk,
	pio_0_external_connection_export);	

	input		clk_clk;
	output	[7:0]	pio_0_external_connection_export;
endmodule
